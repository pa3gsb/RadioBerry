
`include "timescale.v"

module spi_slave(spi_sck, spi_mosi, spi_miso, spi_ce0);


input spi_sck;
input spi_mosi; 
output spi_miso; 
input spi_ce0;






endmodule